module ALU(
  data1_i,
  data2_i,
  ALUCtrl_i,
  data_o,
  Zero_o
);

input signed      [31:0] data1_i;
input signed      [31:0] data2_i;
input              [2:0] ALUCtrl_i;
output reg        [31:0] data_o;
output                   Zero_o; // abandon since not used

`define AND 3'b000
`define XOR 3'b001
`define SLL 3'b010
`define ADD 3'b011
`define SUB 3'b100
`define MUL 3'b101
`define SRAI 3'b110

always@ (*) begin
  case (ALUCtrl_i)
    `AND: data_o <= data1_i & data2_i; 
    `XOR: data_o <= data1_i ^ data2_i;
    `SLL: data_o <= data1_i << data2_i;
    `ADD: data_o <= data1_i + data2_i;
    `SUB: data_o <= data1_i - data2_i;
    `MUL: data_o <= data1_i * data2_i;
    `SRAI: data_o <= data1_i >>> data2_i[4:0];
  endcase
end

endmodule
